`timescale 1 ns/1 ps

module testbench4 ();

reg r_A;
reg r_B;
wire r_Cout;
wire w_S;
wire r_Cin;

endmodule




